Beispil
